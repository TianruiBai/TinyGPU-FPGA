`ifndef UTAH_TEAPOT_DATA_SVH
`define UTAH_TEAPOT_DATA_SVH

// Utah teapot control points and patches (derived from freeglut teapot data, MIT license).
localparam int TEA_INPUT_PATCHES = 10;
localparam int TEA_CP_COUNT = 129;
localparam int teapot_patch [0:TEA_INPUT_PATCHES-1][0:15] = '{
    '{ 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15 },
    '{ 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27 },
    '{ 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 38, 39 },
    '{ 40, 41, 42, 40, 43, 44, 45, 46, 47, 47, 47, 47, 48, 49, 50, 51 },
    '{ 48, 49, 50, 51, 52, 53, 54, 55, 56, 57, 58, 59, 60, 61, 62, 63 },
    '{ 64, 64, 64, 64, 65, 66, 67, 68, 69, 70, 71, 72, 39, 38, 37, 36 },
    '{ 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88 },
    '{ 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100 },
    '{ 101, 102, 103, 104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116 },
    '{ 113, 114, 115, 116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128 }
};

localparam real teapot_cp [0:TEA_CP_COUNT-1][0:2] = '{
    '{ 1.40000, 0.00000, 2.40000 },
    '{ 1.40000, -0.78400, 2.40000 },
    '{ 0.78400, -1.40000, 2.40000 },
    '{ 0.00000, -1.40000, 2.40000 },
    '{ 1.33750, 0.00000, 2.53125 },
    '{ 1.33750, -0.74900, 2.53125 },
    '{ 0.74900, -1.33750, 2.53125 },
    '{ 0.00000, -1.33750, 2.53125 },
    '{ 1.43750, 0.00000, 2.53125 },
    '{ 1.43750, -0.80500, 2.53125 },
    '{ 0.80500, -1.43750, 2.53125 },
    '{ 0.00000, -1.43750, 2.53125 },
    '{ 1.50000, 0.00000, 2.40000 },
    '{ 1.50000, -0.84000, 2.40000 },
    '{ 0.84000, -1.50000, 2.40000 },
    '{ 0.00000, -1.50000, 2.40000 },
    '{ 1.75000, 0.00000, 1.87500 },
    '{ 1.75000, -0.98000, 1.87500 },
    '{ 0.98000, -1.75000, 1.87500 },
    '{ 0.00000, -1.75000, 1.87500 },
    '{ 2.00000, 0.00000, 1.35000 },
    '{ 2.00000, -1.12000, 1.35000 },
    '{ 1.12000, -2.00000, 1.35000 },
    '{ 0.00000, -2.00000, 1.35000 },
    '{ 2.00000, 0.00000, 0.90000 },
    '{ 2.00000, -1.12000, 0.90000 },
    '{ 1.12000, -2.00000, 0.90000 },
    '{ 0.00000, -2.00000, 0.90000 },
    '{ 2.00000, 0.00000, 0.45000 },
    '{ 2.00000, -1.12000, 0.45000 },
    '{ 1.12000, -2.00000, 0.45000 },
    '{ 0.00000, -2.00000, 0.45000 },
    '{ 1.50000, 0.00000, 0.22500 },
    '{ 1.50000, -0.84000, 0.22500 },
    '{ 0.84000, -1.50000, 0.22500 },
    '{ 0.00000, -1.50000, 0.22500 },
    '{ 1.50000, 0.00000, 0.15000 },
    '{ 1.50000, -0.84000, 0.15000 },
    '{ 0.84000, -1.50000, 0.15000 },
    '{ 0.00000, -1.50000, 0.15000 },
    '{ 0.00000, 0.00000, 3.15000 },
    '{ 0.00000, -0.00200, 3.15000 },
    '{ 0.00200, 0.00000, 3.15000 },
    '{ 0.80000, 0.00000, 3.15000 },
    '{ 0.80000, -0.45000, 3.15000 },
    '{ 0.45000, -0.80000, 3.15000 },
    '{ 0.00000, -0.80000, 3.15000 },
    '{ 0.00000, 0.00000, 2.85000 },
    '{ 0.20000, 0.00000, 2.70000 },
    '{ 0.20000, -0.11200, 2.70000 },
    '{ 0.11200, -0.20000, 2.70000 },
    '{ 0.00000, -0.20000, 2.70000 },
    '{ 0.40000, 0.00000, 2.55000 },
    '{ 0.40000, -0.22400, 2.55000 },
    '{ 0.22400, -0.40000, 2.55000 },
    '{ 0.00000, -0.40000, 2.55000 },
    '{ 1.30000, 0.00000, 2.55000 },
    '{ 1.30000, -0.72800, 2.55000 },
    '{ 0.72800, -1.30000, 2.55000 },
    '{ 0.00000, -1.30000, 2.55000 },
    '{ 1.30000, 0.00000, 2.40000 },
    '{ 1.30000, -0.72800, 2.40000 },
    '{ 0.72800, -1.30000, 2.40000 },
    '{ 0.00000, -1.30000, 2.40000 },
    '{ 0.00000, 0.00000, 0.00000 },
    '{ 0.00000, -1.42500, 0.00000 },
    '{ 0.79800, -1.42500, 0.00000 },
    '{ 1.42500, -0.79800, 0.00000 },
    '{ 1.42500, 0.00000, 0.00000 },
    '{ 0.00000, -1.50000, 0.07500 },
    '{ 0.84000, -1.50000, 0.07500 },
    '{ 1.50000, -0.84000, 0.07500 },
    '{ 1.50000, 0.00000, 0.07500 },
    '{ -1.60000, 0.00000, 2.02500 },
    '{ -1.60000, -0.30000, 2.02500 },
    '{ -1.50000, -0.30000, 2.25000 },
    '{ -1.50000, 0.00000, 2.25000 },
    '{ -2.30000, 0.00000, 2.02500 },
    '{ -2.30000, -0.30000, 2.02500 },
    '{ -2.50000, -0.30000, 2.25000 },
    '{ -2.50000, 0.00000, 2.25000 },
    '{ -2.70000, 0.00000, 2.02500 },
    '{ -2.70000, -0.30000, 2.02500 },
    '{ -3.00000, -0.30000, 2.25000 },
    '{ -3.00000, 0.00000, 2.25000 },
    '{ -2.70000, 0.00000, 1.80000 },
    '{ -2.70000, -0.30000, 1.80000 },
    '{ -3.00000, -0.30000, 1.80000 },
    '{ -3.00000, 0.00000, 1.80000 },
    '{ -2.70000, 0.00000, 1.57500 },
    '{ -2.70000, -0.30000, 1.57500 },
    '{ -3.00000, -0.30000, 1.35000 },
    '{ -3.00000, 0.00000, 1.35000 },
    '{ -2.50000, 0.00000, 1.12500 },
    '{ -2.50000, -0.30000, 1.12500 },
    '{ -2.65000, -0.30000, 0.93750 },
    '{ -2.65000, 0.00000, 0.93750 },
    '{ -2.00000, 0.00000, 0.90000 },
    '{ -2.00000, -0.30000, 0.90000 },
    '{ -1.90000, -0.30000, 0.60000 },
    '{ -1.90000, 0.00000, 0.60000 },
    '{ 1.70000, 0.00000, 1.42500 },
    '{ 1.70000, -0.66000, 1.42500 },
    '{ 1.70000, -0.66000, 0.60000 },
    '{ 1.70000, 0.00000, 0.60000 },
    '{ 2.60000, 0.00000, 1.42500 },
    '{ 2.60000, -0.66000, 1.42500 },
    '{ 3.10000, -0.66000, 0.82500 },
    '{ 3.10000, 0.00000, 0.82500 },
    '{ 2.30000, 0.00000, 2.10000 },
    '{ 2.30000, -0.25000, 2.10000 },
    '{ 2.40000, -0.25000, 2.02500 },
    '{ 2.40000, 0.00000, 2.02500 },
    '{ 2.70000, 0.00000, 2.40000 },
    '{ 2.70000, -0.25000, 2.40000 },
    '{ 3.30000, -0.25000, 2.40000 },
    '{ 3.30000, 0.00000, 2.40000 },
    '{ 2.80000, 0.00000, 2.47500 },
    '{ 2.80000, -0.25000, 2.47500 },
    '{ 3.52500, -0.25000, 2.49375 },
    '{ 3.52500, 0.00000, 2.49375 },
    '{ 2.90000, 0.00000, 2.47500 },
    '{ 2.90000, -0.15000, 2.47500 },
    '{ 3.45000, -0.15000, 2.51250 },
    '{ 3.45000, 0.00000, 2.51250 },
    '{ 2.80000, 0.00000, 2.40000 },
    '{ 2.80000, -0.15000, 2.40000 },
    '{ 3.20000, -0.15000, 2.40000 },
    '{ 3.20000, 0.00000, 2.40000 }
};

`endif
