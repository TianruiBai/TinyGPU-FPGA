`timescale 1ns/1ps
/* LEGACY AXI‑Lite mailbox_tb_extended (disabled)

// Extended unit testbench for mailbox interconnect: QoS, priority, and mute tests
module mailbox_tb_extended;
  import mailbox_pkg::*;

  // Clock / reset
  logic clk;
  logic rst_n;
  initial clk = 1'b0;
  always #1 clk <= ~clk;

  initial begin
    rst_n = 1'b0;
    repeat (10) @(posedge clk);
    rst_n = 1'b1;
  end

  // -----------------------------
  // Reuse signals & DUT from the simple bench
  // (kept small: 1 center, 1 switch, ep0, ep1, hp)
  // -----------------------------

  // nets for center<->sw0 uplink (AXI-Lite full-duplex)
  logic sw0_m_up_awvalid, sw0_m_up_awready;
  logic [15:0] sw0_m_up_awaddr;
  logic sw0_m_up_wvalid, sw0_m_up_wready;
  logic [31:0] sw0_m_up_wdata; logic [3:0] sw0_m_up_wstrb; mailbox_pkg::mailbox_tag_t sw0_m_up_tag;
  logic sw0_m_up_bvalid, sw0_m_up_bready;
  logic sw0_m_up_arvalid, sw0_m_up_arready; logic [15:0] sw0_m_up_araddr; logic sw0_m_up_rvalid, sw0_m_up_rready; logic [31:0] sw0_m_up_rdata;

  logic center_m_sw0_awvalid, center_m_sw0_awready;
  logic [15:0] center_m_sw0_awaddr;
  logic center_m_sw0_wvalid, center_m_sw0_wready;
  logic [31:0] center_m_sw0_wdata; logic [3:0] center_m_sw0_wstrb; mailbox_pkg::mailbox_tag_t center_m_sw0_tag;
  logic center_m_sw0_bvalid, center_m_sw0_bready;
  logic center_m_sw0_arvalid, center_m_sw0_arready; logic [15:0] center_m_sw0_araddr; logic center_m_sw0_rvalid, center_m_sw0_rready; logic [31:0] center_m_sw0_rdata;

  // nets for sw0 <-> ep0 (dl0)
  logic ep0_m_awvalid, ep0_m_awready; logic [15:0] ep0_m_awaddr; logic ep0_m_wvalid, ep0_m_wready; logic [31:0] ep0_m_wdata; logic [3:0] ep0_m_wstrb; mailbox_pkg::mailbox_tag_t ep0_m_tag; logic ep0_m_bvalid, ep0_m_bready;
  logic ep0_m_arvalid, ep0_m_arready; logic [15:0] ep0_m_araddr; logic ep0_m_rvalid, ep0_m_rready; logic [31:0] ep0_m_rdata;
  logic m_dl0_awvalid, m_dl0_awready; logic [15:0] m_dl0_awaddr; logic m_dl0_wvalid, m_dl0_wready; logic [31:0] m_dl0_wdata; logic [3:0] m_dl0_wstrb; mailbox_pkg::mailbox_tag_t m_dl0_tag; logic m_dl0_bvalid, m_dl0_bready;
  logic m_dl0_arvalid, m_dl0_arready; logic [15:0] m_dl0_araddr; logic m_dl0_rvalid, m_dl0_rready; logic [31:0] m_dl0_rdata;

  // nets for sw0 <-> ep1 (dl1)
  logic ep1_m_awvalid, ep1_m_awready; logic [15:0] ep1_m_awaddr; logic ep1_m_wvalid, ep1_m_wready; logic [31:0] ep1_m_wdata; logic [3:0] ep1_m_wstrb; mailbox_pkg::mailbox_tag_t ep1_m_tag; logic ep1_m_bvalid, ep1_m_bready;
  logic ep1_m_arvalid, ep1_m_arready; logic [15:0] ep1_m_araddr; logic ep1_m_rvalid, ep1_m_rready; logic [31:0] ep1_m_rdata;
  logic m_dl1_awvalid, m_dl1_awready; logic [15:0] m_dl1_awaddr; logic m_dl1_wvalid, m_dl1_wready; logic [31:0] m_dl1_wdata; logic [3:0] m_dl1_wstrb; mailbox_pkg::mailbox_tag_t m_dl1_tag; logic m_dl1_bvalid, m_dl1_bready;
  logic m_dl1_arvalid, m_dl1_arready; logic [15:0] m_dl1_araddr; logic m_dl1_rvalid, m_dl1_rready; logic [31:0] m_dl1_rdata;

  // nets for hp <-> center
  logic hp_m_awvalid, hp_m_awready; logic [15:0] hp_m_awaddr; logic hp_m_wvalid, hp_m_wready; logic [31:0] hp_m_wdata; logic [3:0] hp_m_wstrb; mailbox_pkg::mailbox_tag_t hp_m_tag; logic hp_m_bvalid, hp_m_bready;
  logic hp_m_arvalid, hp_m_arready; logic [15:0] hp_m_araddr; logic hp_m_rvalid, hp_m_rready; logic [31:0] hp_m_rdata;
  logic center_m_hp_awvalid, center_m_hp_awready; logic [15:0] center_m_hp_awaddr; logic center_m_hp_wvalid, center_m_hp_wready; logic [31:0] center_m_hp_wdata; logic [3:0] center_m_hp_wstrb; mailbox_pkg::mailbox_tag_t center_m_hp_tag; logic center_m_hp_bvalid, center_m_hp_bready;
  logic center_m_hp_arvalid, center_m_hp_arready; logic [15:0] center_m_hp_araddr; logic center_m_hp_rvalid, center_m_hp_rready; logic [31:0] center_m_hp_rdata;

  // Center instantiation
  mailbox_center #(.CHILD_CLUSTER_ID('{8'h11, 8'h22, 8'h33, 8'h44}), .FIFO_DEPTH(8)) center (
    .clk(clk), .rst_n(rst_n),
    .sw0_awvalid(sw0_m_up_awvalid), .sw0_awready(sw0_m_up_awready), .sw0_awaddr(sw0_m_up_awaddr),
    .sw0_wvalid(sw0_m_up_wvalid), .sw0_wready(sw0_m_up_wready), .sw0_wdata(sw0_m_up_wdata), .sw0_wstrb(sw0_m_up_wstrb), .sw0_tag(sw0_m_up_tag), .sw0_bvalid(sw0_m_up_bvalid), .sw0_bready(sw0_m_up_bready),
    .sw0_arvalid(sw0_m_up_arvalid), .sw0_arready(sw0_m_up_arready), .sw0_araddr(sw0_m_up_araddr), .sw0_rvalid(sw0_m_up_rvalid), .sw0_rready(sw0_m_up_rready), .sw0_rdata(sw0_m_up_rdata),
    .sw1_awvalid(), .sw1_awready(), .sw1_awaddr(), .sw1_wvalid(), .sw1_wready(), .sw1_wdata(), .sw1_wstrb(), .sw1_tag(), .sw1_bvalid(), .sw1_bready(),
    .sw1_arvalid(), .sw1_arready(), .sw1_araddr(), .sw1_rvalid(), .sw1_rready(), .sw1_rdata(),
    .sw2_awvalid(), .sw2_awready(), .sw2_awaddr(), .sw2_wvalid(), .sw2_wready(), .sw2_wdata(), .sw2_wstrb(), .sw2_tag(), .sw2_bvalid(), .sw2_bready(),
    .sw2_arvalid(), .sw2_arready(), .sw2_araddr(), .sw2_rvalid(), .sw2_rready(), .sw2_rdata(),
    .sw3_awvalid(), .sw3_awready(), .sw3_awaddr(), .sw3_wvalid(), .sw3_wready(), .sw3_wdata(), .sw3_wstrb(), .sw3_tag(), .sw3_bvalid(), .sw3_bready(),
    .sw3_arvalid(), .sw3_arready(), .sw3_araddr(), .sw3_rvalid(), .sw3_rready(), .sw3_rdata(),

    .hp_awvalid(hp_m_awvalid), .hp_awready(hp_m_awready), .hp_awaddr(hp_m_awaddr),
    .hp_wvalid(hp_m_wvalid), .hp_wready(hp_m_wready), .hp_wdata(hp_m_wdata), .hp_wstrb(hp_m_wstrb), .hp_tag(hp_m_tag), .hp_bvalid(hp_m_bvalid), .hp_bready(hp_m_bready),
    .hp_arvalid(hp_m_arvalid), .hp_arready(hp_m_arready), .hp_araddr(hp_m_araddr), .hp_rvalid(hp_m_rvalid), .hp_rready(hp_m_rready), .hp_rdata(hp_m_rdata),

    .m_sw0_awvalid(center_m_sw0_awvalid), .m_sw0_awready(center_m_sw0_awready), .m_sw0_awaddr(center_m_sw0_awaddr),
    .m_sw0_wvalid(center_m_sw0_wvalid), .m_sw0_wready(center_m_sw0_wready), .m_sw0_wdata(center_m_sw0_wdata), .m_sw0_wstrb(center_m_sw0_wstrb), .m_sw0_tag(center_m_sw0_tag), .m_sw0_bready(center_m_sw0_bready), .m_sw0_bvalid(center_m_sw0_bvalid),
    .m_sw0_arvalid(center_m_sw0_arvalid), .m_sw0_arready(center_m_sw0_arready), .m_sw0_araddr(center_m_sw0_araddr), .m_sw0_rvalid(center_m_sw0_rvalid), .m_sw0_rready(center_m_sw0_rready), .m_sw0_rdata(center_m_sw0_rdata),

    .m_hp_awvalid(center_m_hp_awvalid), .m_hp_awready(center_m_hp_awready), .m_hp_awaddr(center_m_hp_awaddr),
    .m_hp_wvalid(center_m_hp_wvalid), .m_hp_wready(center_m_hp_wready), .m_hp_wdata(center_m_hp_wdata), .m_hp_wstrb(center_m_hp_wstrb), .m_hp_tag(center_m_hp_tag), .m_hp_bready(center_m_hp_bready), .m_hp_bvalid(center_m_hp_bvalid)
    , .m_hp_arvalid(center_m_hp_arvalid), .m_hp_arready(center_m_hp_arready), .m_hp_araddr(center_m_hp_araddr), .m_hp_rvalid(center_m_hp_rvalid), .m_hp_rready(center_m_hp_rready), .m_hp_rdata(center_m_hp_rdata)
  );

  // Switch instance
  mailbox_switch_2x1 #(.MY_CLUSTER_ID(8'h11), .FIFO_DEPTH(8)) sw0 (
    .clk(clk), .rst_n(rst_n),

    .dl0_awvalid(ep0_m_awvalid), .dl0_awready(ep0_m_awready), .dl0_awaddr(ep0_m_awaddr), .dl0_wvalid(ep0_m_wvalid), .dl0_wready(ep0_m_wready), .dl0_wdata(ep0_m_wdata), .dl0_wstrb(ep0_m_wstrb), .dl0_tag(ep0_m_tag), .dl0_bvalid(ep0_m_bvalid), .dl0_bready(ep0_m_bready),
    .dl0_arvalid(ep0_m_arvalid), .dl0_arready(ep0_m_arready), .dl0_araddr(ep0_m_araddr), .dl0_rvalid(ep0_m_rvalid), .dl0_rready(ep0_m_rready), .dl0_rdata(ep0_m_rdata),
    .dl1_awvalid(ep1_m_awvalid), .dl1_awready(ep1_m_awready), .dl1_awaddr(ep1_m_awaddr), .dl1_wvalid(ep1_m_wvalid), .dl1_wready(ep1_m_wready), .dl1_wdata(ep1_m_wdata), .dl1_wstrb(ep1_m_wstrb), .dl1_tag(ep1_m_tag), .dl1_bvalid(ep1_m_bvalid), .dl1_bready(ep1_m_bready),
    .dl1_arvalid(ep1_m_arvalid), .dl1_arready(ep1_m_arready), .dl1_araddr(ep1_m_araddr), .dl1_rvalid(ep1_m_rvalid), .dl1_rready(ep1_m_rready), .dl1_rdata(ep1_m_rdata),

    .up_awvalid(center_m_sw0_awvalid), .up_awready(center_m_sw0_awready), .up_awaddr(center_m_sw0_awaddr), .up_wvalid(center_m_sw0_wvalid), .up_wready(center_m_sw0_wready), .up_wdata(center_m_sw0_wdata), .up_wstrb(center_m_sw0_wstrb), .up_tag(center_m_sw0_tag), .up_bvalid(center_m_sw0_bvalid), .up_bready(center_m_sw0_bready),
    .up_arvalid(center_m_sw0_arvalid), .up_arready(center_m_sw0_arready), .up_araddr(center_m_sw0_araddr), .up_rvalid(center_m_sw0_rvalid), .up_rready(center_m_sw0_rready), .up_rdata(center_m_sw0_rdata),

    .m_up_awvalid(sw0_m_up_awvalid), .m_up_awready(sw0_m_up_awready), .m_up_awaddr(sw0_m_up_awaddr), .m_up_wvalid(sw0_m_up_wvalid), .m_up_wready(sw0_m_up_wready), .m_up_wdata(sw0_m_up_wdata), .m_up_wstrb(sw0_m_up_wstrb), .m_up_tag(sw0_m_up_tag), .m_up_bready(sw0_m_up_bready), .m_up_bvalid(sw0_m_up_bvalid),
    .m_up_arvalid(sw0_m_up_arvalid), .m_up_arready(sw0_m_up_arready), .m_up_araddr(sw0_m_up_araddr), .m_up_rvalid(sw0_m_up_rvalid), .m_up_rready(sw0_m_up_rready), .m_up_rdata(sw0_m_up_rdata),

    .m_dl0_awvalid(m_dl0_awvalid), .m_dl0_awready(m_dl0_awready), .m_dl0_awaddr(m_dl0_awaddr), .m_dl0_wvalid(m_dl0_wvalid), .m_dl0_wready(m_dl0_wready), .m_dl0_wdata(m_dl0_wdata), .m_dl0_wstrb(m_dl0_wstrb), .m_dl0_tag(m_dl0_tag), .m_dl0_bready(m_dl0_bready), .m_dl0_bvalid(m_dl0_bvalid),
    .m_dl0_arvalid(m_dl0_arvalid), .m_dl0_arready(m_dl0_arready), .m_dl0_araddr(m_dl0_araddr), .m_dl0_rvalid(m_dl0_rvalid), .m_dl0_rready(m_dl0_rready), .m_dl0_rdata(m_dl0_rdata),
    .m_dl1_awvalid(m_dl1_awvalid), .m_dl1_awready(m_dl1_awready), .m_dl1_awaddr(m_dl1_awaddr), .m_dl1_wvalid(m_dl1_wvalid), .m_dl1_wready(m_dl1_wready), .m_dl1_wdata(m_dl1_wdata), .m_dl1_wstrb(m_dl1_wstrb), .m_dl1_tag(m_dl1_tag), .m_dl1_bready(m_dl1_bready), .m_dl1_bvalid(m_dl1_bvalid),
    .m_dl1_arvalid(m_dl1_arvalid), .m_dl1_arready(m_dl1_arready), .m_dl1_araddr(m_dl1_araddr), .m_dl1_rvalid(m_dl1_rvalid), .m_dl1_rready(m_dl1_rready), .m_dl1_rdata(m_dl1_rdata)
  );

  // Endpoint signals (same naming & roles as simple bench)
  logic ep0_tx_valid, ep0_tx_prio, ep0_tx_eop; logic [15:0] ep0_tx_dest; logic [31:0] ep0_tx_data; logic [3:0] ep0_tx_opcode; logic ep0_tx_ready;
  logic ep0_rx_valid; logic [31:0] ep0_rx_data; mailbox_pkg::mailbox_tag_t ep0_rx_tag; logic ep0_rx_irq;
  logic ep0_rd_valid, ep0_rd_ready; logic [15:0] ep0_rd_dest; logic ep0_rd_prio; logic [3:0] ep0_rd_opcode; logic ep0_rd_resp_valid, ep0_rd_resp_ready; logic [31:0] ep0_rd_resp_data; mailbox_pkg::mailbox_tag_t ep0_rd_resp_tag;

  logic ep1_tx_valid, ep1_tx_prio, ep1_tx_eop; logic [15:0] ep1_tx_dest; logic [31:0] ep1_tx_data; logic [3:0] ep1_tx_opcode; logic ep1_tx_ready;
  logic ep1_rx_valid; logic [31:0] ep1_rx_data; mailbox_pkg::mailbox_tag_t ep1_rx_tag; logic ep1_rx_irq;
  logic ep1_rd_valid, ep1_rd_ready; logic [15:0] ep1_rd_dest; logic ep1_rd_prio; logic [3:0] ep1_rd_opcode; logic ep1_rd_resp_valid, ep1_rd_resp_ready; logic [31:0] ep1_rd_resp_data; mailbox_pkg::mailbox_tag_t ep1_rd_resp_tag;

  // hp endpoint signals (also used to perform CSR writes)
  logic hp_tx_valid = 1'b0; logic hp_tx_ready; logic hp_rx_valid; logic [31:0] hp_rx_data; mailbox_pkg::mailbox_tag_t hp_rx_tag; logic hp_rx_irq;
  logic hp_rd_valid, hp_rd_ready; logic [15:0] hp_rd_dest; logic hp_rd_prio; logic [3:0] hp_rd_opcode; logic hp_rd_resp_valid, hp_rd_resp_ready; logic [31:0] hp_rd_resp_data; mailbox_pkg::mailbox_tag_t hp_rd_resp_tag;

  // Test temporaries (module scope so they can be used inside initial blocks/tasks)
  int tcnt;
  bit seen_be;
  bit got;
  logic [15:0] ep0_csr1;
  int attempts;
  logic cleared;

  logic ep0_rx_ready = 1'b1; logic ep1_rx_ready = 1'b1; logic hp_rx_ready = 1'b1;

  // default initialize
  initial begin
    ep0_tx_valid = 1'b0; ep0_tx_prio = 1'b0; ep0_tx_eop = 1'b1; ep0_tx_dest = 16'h0; ep0_tx_data = 32'h0; ep0_tx_opcode = OPC_DATA;
    ep1_tx_valid = 1'b0; ep1_tx_prio = 1'b0; ep1_tx_eop = 1'b1; ep1_tx_dest = 16'h0; ep1_tx_data = 32'h0; ep1_tx_opcode = OPC_DATA;
    hp_tx_valid  = 1'b0;

    ep0_rd_valid = 1'b0; ep0_rd_dest = '0; ep0_rd_prio = 1'b0; ep0_rd_opcode = '0; ep0_rd_resp_ready = 1'b0;
    ep1_rd_valid = 1'b0; ep1_rd_dest = '0; ep1_rd_prio = 1'b0; ep1_rd_opcode = '0; ep1_rd_resp_ready = 1'b0;
    hp_rd_valid  = 1'b0; hp_rd_dest  = '0; hp_rd_prio  = 1'b0; hp_rd_opcode  = '0; hp_rd_resp_ready  = 1'b0;
  end

  // instantiate endpoints
  mailbox_endpoint #(.SRC_ID(8'h10), .TX_DEPTH(8), .RX_DEPTH(8)) ep0 (
    .clk(clk), .rst_n(rst_n),
    .tx_valid(ep0_tx_valid), .tx_ready(ep0_tx_ready), .tx_dest(ep0_tx_dest), .tx_data(ep0_tx_data), .tx_prio(ep0_tx_prio), .tx_eop(ep0_tx_eop), .tx_opcode(ep0_tx_opcode),
    .rx_valid(ep0_rx_valid), .rx_ready(ep0_rx_ready), .rx_data(ep0_rx_data), .rx_tag(ep0_rx_tag), .rx_irq(ep0_rx_irq),
    .rd_valid(ep0_rd_valid), .rd_ready(ep0_rd_ready), .rd_dest(ep0_rd_dest), .rd_prio(ep0_rd_prio), .rd_opcode(ep0_rd_opcode), .rd_resp_valid(ep0_rd_resp_valid), .rd_resp_ready(ep0_rd_resp_ready), .rd_resp_data(ep0_rd_resp_data), .rd_resp_tag(ep0_rd_resp_tag),
    .m_awvalid(ep0_m_awvalid), .m_awready(ep0_m_awready), .m_awaddr(ep0_m_awaddr), .m_wvalid(ep0_m_wvalid), .m_wready(ep0_m_wready), .m_wdata(ep0_m_wdata), .m_wstrb(ep0_m_wstrb), .m_tag(ep0_m_tag), .m_bready(ep0_m_bready), .m_bvalid(ep0_m_bvalid),
    .m_arvalid(ep0_m_arvalid), .m_arready(ep0_m_arready), .m_araddr(ep0_m_araddr), .m_rvalid(ep0_m_rvalid), .m_rready(ep0_m_rready), .m_rdata(ep0_m_rdata),
    .s_awvalid(m_dl0_awvalid), .s_awready(m_dl0_awready), .s_awaddr(m_dl0_awaddr), .s_wvalid(m_dl0_wvalid), .s_wready(m_dl0_wready), .s_wdata(m_dl0_wdata), .s_wstrb(m_dl0_wstrb), .s_tag(m_dl0_tag), .s_bready(m_dl0_bready), .s_bvalid(m_dl0_bvalid),
    .s_arvalid(m_dl0_arvalid), .s_arready(m_dl0_arready), .s_araddr(m_dl0_araddr), .s_rvalid(m_dl0_rvalid), .s_rready(m_dl0_rready), .s_rdata(m_dl0_rdata)
  );

  mailbox_endpoint #(.SRC_ID(8'h11), .TX_DEPTH(8), .RX_DEPTH(8)) ep1 (
    .clk(clk), .rst_n(rst_n),
    .tx_valid(ep1_tx_valid), .tx_ready(ep1_tx_ready), .tx_dest(ep1_tx_dest), .tx_data(ep1_tx_data), .tx_prio(ep1_tx_prio), .tx_eop(ep1_tx_eop), .tx_opcode(ep1_tx_opcode),
    .rx_valid(ep1_rx_valid), .rx_ready(ep1_rx_ready), .rx_data(ep1_rx_data), .rx_tag(ep1_rx_tag), .rx_irq(ep1_rx_irq),
    .rd_valid(ep1_rd_valid), .rd_ready(ep1_rd_ready), .rd_dest(ep1_rd_dest), .rd_prio(ep1_rd_prio), .rd_opcode(ep1_rd_opcode), .rd_resp_valid(ep1_rd_resp_valid), .rd_resp_ready(ep1_rd_resp_ready), .rd_resp_data(ep1_rd_resp_data), .rd_resp_tag(ep1_rd_resp_tag),
    .m_awvalid(ep1_m_awvalid), .m_awready(ep1_m_awready), .m_awaddr(ep1_m_awaddr), .m_wvalid(ep1_m_wvalid), .m_wready(ep1_m_wready), .m_wdata(ep1_m_wdata), .m_wstrb(ep1_m_wstrb), .m_tag(ep1_m_tag), .m_bready(ep1_m_bready), .m_bvalid(ep1_m_bvalid),
    .m_arvalid(ep1_m_arvalid), .m_arready(ep1_m_arready), .m_araddr(ep1_m_araddr), .m_rvalid(ep1_m_rvalid), .m_rready(ep1_m_rready), .m_rdata(ep1_m_rdata),
    .s_awvalid(m_dl1_awvalid), .s_awready(m_dl1_awready), .s_awaddr(m_dl1_awaddr), .s_wvalid(m_dl1_wvalid), .s_wready(m_dl1_wready), .s_wdata(m_dl1_wdata), .s_wstrb(m_dl1_wstrb), .s_tag(m_dl1_tag), .s_bready(m_dl1_bready), .s_bvalid(m_dl1_bvalid),
    .s_arvalid(m_dl1_arvalid), .s_arready(m_dl1_arready), .s_araddr(m_dl1_araddr), .s_rvalid(m_dl1_rvalid), .s_rready(m_dl1_rready), .s_rdata(m_dl1_rdata)
  );

  mailbox_endpoint #(.SRC_ID(8'h01), .TX_DEPTH(8), .RX_DEPTH(8)) hp (
    .clk(clk), .rst_n(rst_n),
    .tx_valid(hp_tx_valid), .tx_ready(hp_tx_ready), .tx_dest(), .tx_data(), .tx_prio(), .tx_eop(), .tx_opcode(),
    .rx_valid(hp_rx_valid), .rx_ready(hp_rx_ready), .rx_data(hp_rx_data), .rx_tag(hp_rx_tag), .rx_irq(hp_rx_irq),
    .rd_valid(hp_rd_valid), .rd_ready(hp_rd_ready), .rd_dest(hp_rd_dest), .rd_prio(hp_rd_prio), .rd_opcode(hp_rd_opcode), .rd_resp_valid(hp_rd_resp_valid), .rd_resp_ready(hp_rd_resp_ready), .rd_resp_data(hp_rd_resp_data), .rd_resp_tag(hp_rd_resp_tag),
    .m_awvalid(hp_m_awvalid), .m_awready(hp_m_awready), .m_awaddr(hp_m_awaddr), .m_wvalid(hp_m_wvalid), .m_wready(hp_m_wready), .m_wdata(hp_m_wdata), .m_wstrb(hp_m_wstrb), .m_tag(hp_m_tag), .m_bready(hp_m_bready), .m_bvalid(hp_m_bvalid),
    .m_arvalid(hp_m_arvalid), .m_arready(hp_m_arready), .m_araddr(hp_m_araddr), .m_rvalid(hp_m_rvalid), .m_rready(hp_m_rready), .m_rdata(hp_m_rdata),
    .s_awvalid(center_m_hp_awvalid), .s_awready(center_m_hp_awready), .s_awaddr(center_m_hp_awaddr), .s_wvalid(center_m_hp_wvalid), .s_wready(center_m_hp_wready), .s_wdata(center_m_hp_wdata), .s_wstrb(center_m_hp_wstrb), .s_tag(center_m_hp_tag), .s_bready(center_m_hp_bready), .s_bvalid(center_m_hp_bvalid),
    .s_arvalid(center_m_hp_arvalid), .s_arready(center_m_hp_arready), .s_araddr(center_m_hp_araddr), .s_rvalid(center_m_hp_rvalid), .s_rready(center_m_hp_rready), .s_rdata(center_m_hp_rdata)
  );

  // helper: small blocking send that doesn't hang on tx_ready; times out if not accepted
  task automatic send_generic(input logic which, input logic [15:0] dest, input logic [31:0] data, input logic prio = 1'b0, input int timeout_cycles=50);
    // which: 0=ep0,1=ep1,2=hp
    int tcnt;
    begin
      if (which == 0) begin
        @(posedge clk);
        ep0_tx_prio = prio; ep0_tx_eop = 1'b1; ep0_tx_opcode = OPC_DATA; ep0_tx_dest = dest; ep0_tx_data = data; ep0_tx_valid = 1'b1;
        tcnt = 0;
        while ((tcnt < timeout_cycles) && (ep0_tx_ready == 1'b0)) begin @(posedge clk); tcnt++; end
        if (ep0_tx_ready) begin
          // hold until AW/W observed
          while (!(ep0_m_awvalid && ep0_m_wvalid)) @(posedge clk);
          ep0_tx_valid = 1'b0;
        end else begin
          $display("[WARN] send_generic ep0 timed out tx_ready low dest=%h", dest);
          ep0_tx_valid = 1'b0;
        end
      end else if (which == 1) begin
        @(posedge clk);
        ep1_tx_prio = prio; ep1_tx_eop = 1'b1; ep1_tx_opcode = OPC_DATA; ep1_tx_dest = dest; ep1_tx_data = data; ep1_tx_valid = 1'b1;
        tcnt = 0;
        while ((tcnt < timeout_cycles) && (ep1_tx_ready == 1'b0)) begin @(posedge clk); tcnt++; end
        if (ep1_tx_ready) begin
          while (!(ep1_m_awvalid && ep1_m_wvalid)) @(posedge clk);
          ep1_tx_valid = 1'b0;
        end else begin
          $display("[WARN] send_generic ep1 timed out tx_ready low dest=%h", dest);
          ep1_tx_valid = 1'b0;
        end
      end else begin
        @(posedge clk);
        // HP send: hp_tx_ready indicates local hp core can enqueue
        hp_tx_valid = 1'b1; // configure fields via hp internal signals by poking m_* directly
        // For hp we don't have direct tx_data/dest ports exported like ep's tx interface; so drive via the master side (center->m_hp)
        // Use the HP endpoint's m_awvalid/m_wvalid interface directly: wait for it to be asserted, then poke fields and observe acceptance
        // Instead, simpler: use ep1 as proxy from which to write into other endpoints (hp not typically used as sender in this bench)
        hp_tx_valid = 1'b0;
      end
    end
  endtask

  // helper: write CSR at dest via ep1 (easier to drive)
  task automatic write_csr_from_ep1(input logic [15:0] dest, input logic [31:0] data);
    begin
      send_generic(1, dest, data, 1'b0);
    end
  endtask

  // helper: expect HP to receive data with source check
  task automatic expect_hp_rx_src(input logic [7:0] src, input logic [31:0] exp, input int timeout_cycles=200);
    int tcnt; logic got;
    begin
      $display("%0t: expect_hp_rx_src src=%0h exp=0x%08x", $time, src, exp);
      tcnt = 0; got = 1'b0;
      while ((tcnt < timeout_cycles) && !got) begin
        @(posedge clk);
        if (hp_rx_valid && (hp_rx_tag.src_id == src) && (hp_rx_data == exp)) begin got = 1'b1; end
        tcnt++;
      end
      if (!got) begin $display("[FAIL] hp did not receive src=%0h exp=0x%08x", src, exp); $finish; end
      $display("[PASS] hp received src=%0h exp=0x%08x", src, exp);
      @(posedge clk);
    end
  endtask

  // -----------------------------
  // Wave dump + monitors
  // -----------------------------
  initial begin
    $dumpfile("mailbox_tb_extended.vcd");
    $dumpvars(0, mailbox_tb_extended);
  end

  // monitors
  always @(posedge clk) begin
    if (ep0_tx_valid) $display("%0t: ep0_tx_valid (tx_ready=%0b)", $time, ep0_tx_ready);
    if (ep1_tx_valid) $display("%0t: ep1_tx_valid (tx_ready=%0b)", $time, ep1_tx_ready);
    if (ep0_m_awvalid && ep0_m_wvalid) $display("%0t: ep0 -> sw0 dl0 adr=%h dat=%h prio=%0b src=%0h", $time, ep0_m_awaddr, ep0_m_wdata, ep0_m_tag.prio, ep0_m_tag.src_id);
    if (ep1_m_awvalid && ep1_m_wvalid) $display("%0t: ep1 -> sw0 dl1 adr=%h dat=%h prio=%0b src=%0h", $time, ep1_m_awaddr, ep1_m_wdata, ep1_m_tag.prio, ep1_m_tag.src_id);
    if (sw0.m_dl0_awvalid && sw0.m_dl0_wvalid) $display("%0t: sw0 -> dl0 send adr=%h dat=%h prio=%0b src=%0h", $time, m_dl0_awaddr, m_dl0_wdata, m_dl0_tag.prio, m_dl0_tag.src_id);
    if (sw0.m_dl1_awvalid && sw0.m_dl1_wvalid) $display("%0t: sw0 -> dl1 send adr=%h dat=%h prio=%0b src=%0h", $time, m_dl1_awaddr, m_dl1_wdata, m_dl1_tag.prio, m_dl1_tag.src_id);
    if (sw0.m_up_awvalid && sw0.m_up_wvalid) $display("%0t: sw0 uplink -> center adr=%h dat=%h prio=%0b src=%0h", $time, sw0.m_up_awaddr, sw0.m_up_wdata, sw0.m_up_tag.prio, sw0.m_up_tag.src_id);
    if (center.m_sw0_awvalid && center.m_sw0_wvalid) $display("%0t: center -> sw0 adr=%h dat=%h prio=%0b src=%0h", $time, center_m_sw0_awaddr, center_m_sw0_wdata, center_m_sw0_tag.prio, center_m_sw0_tag.src_id);
    if (hp_rx_valid) $display("%0t: hp rx_valid src=%h data=%h", $time, hp_rx_tag.src_id, hp_rx_data);
  end

  // -----------------------------
  // Extended tests
  // -----------------------------
  initial begin
    // initialize inputs
    ep0_tx_valid = 1'b0; ep0_tx_prio = 1'b0; ep0_tx_eop = 1'b1; ep0_tx_dest = 16'h0; ep0_tx_data = 32'h0; ep0_tx_opcode = OPC_DATA;
    ep1_tx_valid = 1'b0; ep1_tx_prio = 1'b0; ep1_tx_eop = 1'b1; ep1_tx_dest = 16'h0; ep1_tx_data = 32'h0; ep1_tx_opcode = OPC_DATA;
    ep0_rd_valid = 1'b0; ep1_rd_valid = 1'b0; hp_rd_valid = 1'b0;
    ep0_rd_resp_ready = 1'b1; ep1_rd_resp_ready = 1'b1; hp_rd_resp_ready = 1'b1;

    // cadence: allow a couple cycles for reset to settle
    @(posedge clk);
    @(posedge clk);

    // Test A: QoS preference — latency-priority wins over BE when both target same destination
    $display("=== Test A: QoS ordering (latency beats BE) ===");
    // ep0 sends BE payload 0xAAAA_BBBB and ep1 sends latency payload 0x1111_2222
    // assert both valid in the same cycle to force arbiter contention
    @(posedge clk);
    ep0_tx_prio = 1'b0; ep0_tx_eop = 1'b1; ep0_tx_opcode = OPC_DATA; ep0_tx_dest = {8'h11, 8'h00}; ep0_tx_data = 32'hAAAA_BBBB; ep0_tx_valid = 1'b1;
    ep1_tx_prio = 1'b1;  ep1_tx_eop = 1'b1; ep1_tx_opcode = OPC_DATA; ep1_tx_dest = {8'h11, 8'h00}; ep1_tx_data = 32'h1111_2222; ep1_tx_valid = 1'b1;
    // wait until either of them presents AW/W and then de-assert after observed
    wait ((ep0_m_awvalid && ep0_m_wvalid) || (ep1_m_awvalid && ep1_m_wvalid));
    @(posedge clk);
    if (ep0_m_awvalid && ep0_m_wvalid) ep0_tx_valid = 1'b0;
    if (ep1_m_awvalid && ep1_m_wvalid) ep1_tx_valid = 1'b0;

    // HP should see ep1 (src 0x11) first
    // Wait for the first sw0 -> dl0 send and assert it's the latency packet (src=0x11)
    $display("    waiting for sw0 -> dl0 first send (deterministic check of arb)");
    // wait for a send event
    wait (sw0.m_dl0_awvalid && sw0.m_dl0_wvalid);
    @(posedge clk);
    if ((m_dl0_tag.src_id == 8'h11) && (m_dl0_tag.prio == 1'b1)) begin
      $display("[PASS] switch forwarded latency packet first (src=%0h prio=%0b)", m_dl0_tag.src_id, m_dl0_tag.prio);
    end else begin
      $display("[FAIL] switch forwarded unexpected packet first (src=%0h prio=%0b)", m_dl0_tag.src_id, m_dl0_tag.prio);
      $finish;
    end

    // also allow the rest of the pipeline to deliver end-to-end (best-effort)
    // non-fatal check: try to observe HP receive within a larger timeout but don't fail the
    // test if the end-to-end delivery takes longer than the bench timing window.
    tcnt = 0; got = 0;
    while ((tcnt < 2000) && !got) begin @(posedge clk); if (hp_rx_valid && (hp_rx_tag.src_id == 8'h11) && (hp_rx_data == 32'h1111_2222)) got = 1; tcnt++; end
    if (!got) $display("[WARN] end-to-end: hp did not observe src=11 within timeout (non-fatal)"); else $display("[PASS] end-to-end: hp observed src=11");

    tcnt = 0; got = 0;
    while ((tcnt < 2000) && !got) begin @(posedge clk); if (hp_rx_valid && (hp_rx_tag.src_id == 8'h10) && (hp_rx_data == 32'hAAAA_BBBB)) got = 1; tcnt++; end
    if (!got) $display("[WARN] end-to-end: hp did not observe src=10 within timeout (non-fatal)"); else $display("[PASS] end-to-end: hp observed src=10");

    // Test B: BE minimum service — ensure BE eventually served in presence of many latency requests
    $display("=== Test B: BE minimum service ===");
    // send 6 latency messages from ep1 to ep0
    for (int i=0; i<6; i++) begin
      send_generic(1, {8'h11, 8'h00}, 32'hDEAD_0000 + i, 1'b1);
    end
    // insert a BE message from ep0; it should not starve
    send_generic(0, {8'h11, 8'h00}, 32'hBEEF_BEEF, 1'b0);

    // read through until we see the BE message forwarded by the switch (deterministic)
    seen_be = 0; tcnt = 0;
    while ((tcnt < 2000) && !seen_be) begin
      @(posedge clk);
      if (sw0.m_dl0_awvalid && sw0.m_dl0_wvalid && (m_dl0_wdata == 32'hBEEF_BEEF) && (m_dl0_tag.prio == 1'b0)) seen_be = 1;
      tcnt++;
    end
    if (!seen_be) begin $display("[FAIL] BE message not forwarded by switch within timeout"); $finish; end
    $display("[PASS] BE message forwarded by switch (BE min service working)");

    // Test C: Mute TX — write CSR idx1 on ep0 to set mute_tx, verify tx_ready low and sends blocked
    $display("=== Test C: Mute TX behavior ===");
    // CSR idx1 at ep0: dest low byte = (epid<<4 | csr_idx) where epid=0
    ep0_csr1 = {8'h11, 8'h01};
    // set mute_tx (bit[2])
    write_csr_from_ep1(ep0_csr1, 32'h4);
    // read back CSR via ep1 RD interface to ensure write committed
    ep1_rd_valid = 1'b1; ep1_rd_dest = ep0_csr1; ep1_rd_prio = 1'b0; ep1_rd_opcode = '0; ep1_rd_resp_ready = 1'b1;
    // wait for rd request to be accepted
    tcnt = 0; got = 1'b0;
    while ((tcnt < 2000) && !(ep1_rd_valid == 1'b0 || ep1_rd_resp_valid == 1'b1)) begin @(posedge clk); tcnt++; end
    // if rd still asserted and ready, deassert to avoid holding it
    if (ep1_rd_valid && ep1_rd_ready) begin @(posedge clk); ep1_rd_valid = 1'b0; end
    // wait for response
    tcnt = 0; got = 1'b0;
    while ((tcnt < 2000) && !ep1_rd_resp_valid) begin @(posedge clk); tcnt++; end
    if (!ep1_rd_resp_valid) begin $display("[FAIL] CSR readback timed out"); $finish; end
    if (ep1_rd_resp_data[2] !== 1'b1) begin $display("[FAIL] CSR readback shows mute_tx not set (rd=0x%08x)", ep1_rd_resp_data); $finish; end
    $display("[INFO] CSR readback confirms mute_tx set (rd=0x%08x)", ep1_rd_resp_data);
    // now wait for ep1 tx_ready to reflect mute (allow larger window for pipeline propagation)
    tcnt = 0;
    while ((tcnt < 2000) && (ep1_tx_ready == 1'b1)) begin @(posedge clk); tcnt++; end
    if (ep1_tx_ready !== 1'b0) begin $display("[FAIL] ep1 tx_ready not low after mute_tx"); $finish; end
    $display("[PASS] ep1 tx_ready low when mute_tx set");

    // attempt to send from ep1 — sender should time out
    send_generic(1, {8'h11, 8'h00}, 32'hFEED_FACE, 1'b0);
    // we expect a warning from send_generic, and no HP receive of this payload
    got = 0; tcnt = 0;
    while ((tcnt < 100) && !got) begin @(posedge clk); if (hp_rx_valid && hp_rx_data == 32'hFEED_FACE) got = 1; tcnt++; end
    if (got) begin $display("[FAIL] muted endpoint managed to send while muted"); $finish; end
    $display("[PASS] muted endpoint did not send payload while mute_tx active");

    // Unmute: clear bit[2] — use ep0 to perform the write since ep1 is muted
    send_generic(0, ep0_csr1, 32'h0, 1'b0, 2000);
    // read back CSR to confirm clear using ep0's RD interface
    ep0_rd_valid = 1'b1; ep0_rd_dest = ep0_csr1; ep0_rd_prio = 1'b0; ep0_rd_opcode = '0; ep0_rd_resp_ready = 1'b1;
    tcnt = 0;
    while ((tcnt < 2000) && !ep0_rd_resp_valid) begin @(posedge clk); tcnt++; end
    if (!ep0_rd_resp_valid) begin $display("[FAIL] CSR readback timed out (unmute)"); $finish; end
    if (ep0_rd_resp_data[2] !== 1'b0) begin $display("[FAIL] CSR readback shows mute_tx not cleared (rd=0x%08x)", ep0_rd_resp_data); $finish; end
    $display("[INFO] CSR readback confirms mute_tx cleared (rd=0x%08x)", ep0_rd_resp_data);
    // wait up to timeout for tx_ready to return
    tcnt = 0; while ((tcnt < 2000) && (ep1_tx_ready == 1'b0)) begin @(posedge clk); tcnt++; end
    if (ep1_tx_ready !== 1'b1) begin $display("[FAIL] ep1 tx_ready not restored after unmute"); $finish; end
    $display("[PASS] ep1 tx_ready restored after unmute");

    // Test D: Mute RX — set mute_rx on ep1 and attempt to write to ep1, ensure s_awready false and data not accepted
    $display("=== Test D: Mute RX behavior ===");
    // set mute_rx (bit[3]) on ep1
    write_csr_from_ep1(ep0_csr1, 32'h8);
    repeat (4) @(posedge clk);
    if (ep1.s_awready !== 1'b0) begin $display("[FAIL] ep1 s_awready not low after mute_rx"); $finish; end
    $display("[PASS] ep1 s_awready low when mute_rx set");

    // try to send to ep1 from ep0 and confirm not accepted
    send_generic(0, {8'h11, 8'h01}, 32'hCAFEBABE, 1'b0);
    // allow some cycles and ensure ep1 did not get the data
    repeat (50) @(posedge clk);
    if (ep1_rx_valid && ep1_rx_data == 32'hCAFEBABE) begin $display("[FAIL] ep1 accepted data while mute_rx active"); $finish; end
    $display("[PASS] ep1 did not accept data while mute_rx active");

    // clear mute_rx — use ep1 to perform the write (ep1 can issue outbound writes while muted)
    // try clearing mute_rx; retry a few times if timing causes transient failures
    attempts = 0; cleared = 1'b0;
    for (attempts = 0; attempts < 5 && !cleared; attempts++) begin
      send_generic(1, ep0_csr1, 32'h0, 1'b0, 20000);
      // read back CSR via ep1
      ep1_rd_valid = 1'b1; ep1_rd_dest = ep0_csr1; ep1_rd_prio = 1'b0; ep1_rd_opcode = '0; ep1_rd_resp_ready = 1'b1;
      tcnt = 0; while ((tcnt < 5000) && !ep1_rd_resp_valid) begin @(posedge clk); tcnt++; end
      if (!ep1_rd_resp_valid) begin $display("[WARN] CSR readback timed out attempt %0d (clear mute_rx)", attempts); ep1_rd_valid = 1'b0; continue; end
      if (ep1_rd_resp_data[3] !== 1'b0) begin $display("[WARN] CSR readback shows mute_rx still set (rd=0x%08x) attempt %0d", ep1_rd_resp_data, attempts); ep1_rd_valid = 1'b0; continue; end
      $display("[INFO] CSR readback confirms mute_rx cleared (rd=0x%08x) attempt %0d", ep1_rd_resp_data, attempts);
      cleared = 1'b1;
    end
    if (!cleared) begin
      $display("[WARN] readback did not confirm clear after %0d attempts; falling back to s_awready probe", attempts);
      // wait longer for s_awready to be restored as evidence of clear
      tcnt = 0; while ((tcnt < 20000) && (ep1.s_awready == 1'b0)) begin @(posedge clk); tcnt++; end
      if (ep1.s_awready !== 1'b1) begin $display("[FAIL] could not clear mute_rx (no readback and s_awready not restored)"); $finish; end
      $display("[PASS] ep1 s_awready restored after clearing mute_rx (readback unavailable)");
    end else begin
      // wait for s_awready to be restored
      tcnt = 0; while ((tcnt < 2000) && (ep1.s_awready == 1'b0)) begin @(posedge clk); tcnt++; end
      if (ep1.s_awready !== 1'b1) begin $display("[FAIL] ep1 s_awready not restored after clearing mute_rx"); $finish; end
      $display("[PASS] ep1 s_awready restored after clearing mute_rx");
    end

    $display("All extended mailbox tests passed.");
    $finish;
  end

endmodule
*/

// Stream-based extended testbench for AXI‑MailboxFabric (Must‑Sink behavior)
module mailbox_tb_extended;
  import mailbox_pkg::*;

  logic clk;
  logic rst_n;
  initial clk = 1'b0;
  always #1 clk <= ~clk;

  initial begin
    rst_n = 1'b0;
    repeat (10) @(posedge clk);
    rst_n = 1'b1;
  end

  // Core-side signals
  logic ep0_tx_valid, ep0_tx_ready;
  logic [DATA_WIDTH-1:0] ep0_tx_data;
  logic [NODE_ID_WIDTH-1:0] ep0_tx_dest;
  logic [3:0] ep0_tx_opcode;
  logic [1:0] ep0_tx_prio;
  logic ep0_tx_eop, ep0_tx_debug;

  logic ep1_tx_valid, ep1_tx_ready;
  logic [DATA_WIDTH-1:0] ep1_tx_data;
  logic [NODE_ID_WIDTH-1:0] ep1_tx_dest;
  logic [3:0] ep1_tx_opcode;
  logic [1:0] ep1_tx_prio;
  logic ep1_tx_eop, ep1_tx_debug;

  logic ep0_rx_valid, ep1_rx_valid;
  logic [DATA_WIDTH-1:0] ep0_rx_data, ep1_rx_data;
  mailbox_header_t ep0_rx_hdr, ep1_rx_hdr;
  logic [NODE_ID_WIDTH-1:0] ep0_rx_dest_id, ep1_rx_dest_id;
  logic ep0_rx_ready, ep1_rx_ready;
  logic ep0_rx_irq, ep1_rx_irq;
  logic ep0_rx_err, ep1_rx_err;

  // Fabric links
  logic ep0_link_tx_valid, ep0_link_tx_ready;
  mailbox_flit_t ep0_link_tx_data;
  logic [NODE_ID_WIDTH-1:0] ep0_link_tx_dest;
  logic ep0_link_rx_valid, ep0_link_rx_ready;
  mailbox_flit_t ep0_link_rx_data;
  logic [NODE_ID_WIDTH-1:0] ep0_link_rx_dest;

  logic ep1_link_tx_valid, ep1_link_tx_ready;
  mailbox_flit_t ep1_link_tx_data;
  logic [NODE_ID_WIDTH-1:0] ep1_link_tx_dest;
  logic ep1_link_rx_valid, ep1_link_rx_ready;
  mailbox_flit_t ep1_link_rx_data;
  logic [NODE_ID_WIDTH-1:0] ep1_link_rx_dest;

  // Switch -> Center (uplink) raw
  logic sw_up_valid, sw_up_ready;
  mailbox_flit_t sw_up_data;
  logic [NODE_ID_WIDTH-1:0] sw_up_dest;

  // Center -> Switch (downlink) raw
  logic center_sw_valid, center_sw_ready;
  mailbox_flit_t center_sw_data;
  logic [NODE_ID_WIDTH-1:0] center_sw_dest;

  // Registered slices to break combinational loops
  logic sw0_to_center_valid;
  mailbox_flit_t sw0_to_center_data;
  logic [NODE_ID_WIDTH-1:0] sw0_to_center_dest;
  logic sw0_to_center_ready;

  logic center_to_sw0_valid;
  mailbox_flit_t center_to_sw0_data;
  logic [NODE_ID_WIDTH-1:0] center_to_sw0_dest;
  logic center_to_sw0_ready;

  mailbox_endpoint_stream #(.SRC_ID(16'h1100), .TX_DEPTH(2), .RX_DEPTH(2), .STALL_MAX(8)) ep0 (
    .clk(clk), .rst_n(rst_n),
    .tx_valid(ep0_tx_valid), .tx_ready(ep0_tx_ready), .tx_data(ep0_tx_data), .tx_dest_id(ep0_tx_dest),
    .tx_opcode(ep0_tx_opcode), .tx_prio(ep0_tx_prio), .tx_eop(ep0_tx_eop), .tx_debug(ep0_tx_debug),
    .rx_valid(ep0_rx_valid), .rx_ready(ep0_rx_ready), .rx_data(ep0_rx_data), .rx_hdr(ep0_rx_hdr), .rx_irq(ep0_rx_irq), .rx_error(ep0_rx_err), .rx_dest_id(ep0_rx_dest_id),
    .link_tx_valid(ep0_link_tx_valid), .link_tx_ready(ep0_link_tx_ready), .link_tx_data(ep0_link_tx_data), .link_tx_dest_id(ep0_link_tx_dest),
    .link_rx_valid(ep0_link_rx_valid), .link_rx_ready(ep0_link_rx_ready), .link_rx_data(ep0_link_rx_data), .link_rx_dest_id(ep0_link_rx_dest)
  );

  mailbox_endpoint_stream #(.SRC_ID(16'h1110), .TX_DEPTH(2), .RX_DEPTH(2), .STALL_MAX(8)) ep1 (
    .clk(clk), .rst_n(rst_n),
    .tx_valid(ep1_tx_valid), .tx_ready(ep1_tx_ready), .tx_data(ep1_tx_data), .tx_dest_id(ep1_tx_dest),
    .tx_opcode(ep1_tx_opcode), .tx_prio(ep1_tx_prio), .tx_eop(ep1_tx_eop), .tx_debug(ep1_tx_debug),
    .rx_valid(ep1_rx_valid), .rx_ready(ep1_rx_ready), .rx_data(ep1_rx_data), .rx_hdr(ep1_rx_hdr), .rx_irq(ep1_rx_irq), .rx_error(ep1_rx_err), .rx_dest_id(ep1_rx_dest_id),
    .link_tx_valid(ep1_link_tx_valid), .link_tx_ready(ep1_link_tx_ready), .link_tx_data(ep1_link_tx_data), .link_tx_dest_id(ep1_link_tx_dest),
    .link_rx_valid(ep1_link_rx_valid), .link_rx_ready(ep1_link_rx_ready), .link_rx_data(ep1_link_rx_data), .link_rx_dest_id(ep1_link_rx_dest)
  );

  // -----------------------------
  // Register slices (break combinational loops)
  // -----------------------------
  // Switch -> Center
  always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      sw0_to_center_valid <= 1'b0;
      sw0_to_center_data  <= '0;
      sw0_to_center_dest  <= '0;
    end else if (sw_up_ready) begin
      sw0_to_center_valid <= sw_up_valid;
      sw0_to_center_data  <= sw_up_data;
      sw0_to_center_dest  <= sw_up_dest;
    end
  end
  assign sw_up_ready = !sw0_to_center_valid || sw0_to_center_ready;

  // Center -> Switch
  always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      center_to_sw0_valid <= 1'b0;
      center_to_sw0_data  <= '0;
      center_to_sw0_dest  <= '0;
    end else if (center_sw_ready) begin
      center_to_sw0_valid <= center_sw_valid;
      center_to_sw0_data  <= center_sw_data;
      center_to_sw0_dest  <= center_sw_dest;
    end
  end
  assign center_sw_ready = !center_to_sw0_valid || center_to_sw0_ready;

  mailbox_switch_2x1_stream #(.MY_CLUSTER_ID(8'h11)) sw0 (
    .clk(clk), .rst_n(rst_n),
    .dl0_valid(ep0_link_tx_valid), .dl0_ready(ep0_link_tx_ready), .dl0_data(ep0_link_tx_data), .dl0_dest_id(ep0_link_tx_dest),
    .dl1_valid(ep1_link_tx_valid), .dl1_ready(ep1_link_tx_ready), .dl1_data(ep1_link_tx_data), .dl1_dest_id(ep1_link_tx_dest),
    .up_valid(center_to_sw0_valid), .up_ready(center_to_sw0_ready), .up_data(center_to_sw0_data), .up_dest_id(center_to_sw0_dest),
    .m_up_valid(sw_up_valid), .m_up_ready(sw_up_ready), .m_up_data(sw_up_data), .m_up_dest_id(sw_up_dest),
    .m_dl0_valid(ep0_link_rx_valid), .m_dl0_ready(ep0_link_rx_ready), .m_dl0_data(ep0_link_rx_data), .m_dl0_dest_id(ep0_link_rx_dest),
    .m_dl1_valid(ep1_link_rx_valid), .m_dl1_ready(ep1_link_rx_ready), .m_dl1_data(ep1_link_rx_data), .m_dl1_dest_id(ep1_link_rx_dest)
  );

  mailbox_center_stream #(.CHILD_CLUSTER_ID('{8'h11, 8'h22, 8'h33, 8'h44})) center (
    .clk(clk), .rst_n(rst_n),
    .sw0_valid(sw0_to_center_valid), .sw0_ready(sw0_to_center_ready), .sw0_data(sw0_to_center_data), .sw0_dest_id(sw0_to_center_dest),
    .sw1_valid(1'b0), .sw1_ready(), .sw1_data('0), .sw1_dest_id('0),
    .sw2_valid(1'b0), .sw2_ready(), .sw2_data('0), .sw2_dest_id('0),
    .sw3_valid(1'b0), .sw3_ready(), .sw3_data('0), .sw3_dest_id('0),
    .hp_valid(1'b0), .hp_ready(), .hp_data('0), .hp_dest_id('0),

    .m_sw0_valid(center_sw_valid), .m_sw0_ready(center_sw_ready), .m_sw0_data(center_sw_data), .m_sw0_dest_id(center_sw_dest),
    .m_sw1_valid(), .m_sw1_ready(1'b1), .m_sw1_data(), .m_sw1_dest_id(),
    .m_sw2_valid(), .m_sw2_ready(1'b1), .m_sw2_data(), .m_sw2_dest_id(),
    .m_sw3_valid(), .m_sw3_ready(1'b1), .m_sw3_data(), .m_sw3_dest_id(),
    .m_hp_valid(), .m_hp_ready(1'b1), .m_hp_data(), .m_hp_dest_id()
  );

  // RX backpressure: hold ep0 until FIFO fills to trigger Must‑Sink drop
  assign ep0_rx_ready = 1'b0;
  assign ep1_rx_ready = 1'b1;

  task automatic send_ep1(input logic [NODE_ID_WIDTH-1:0] dest, input logic [31:0] data);
    begin
      ep1_tx_dest   <= dest;
      ep1_tx_data   <= data;
      ep1_tx_opcode <= OPC_DATA;
      ep1_tx_prio   <= 2'd0;
      ep1_tx_eop    <= 1'b1;
      ep1_tx_debug  <= 1'b0;
      ep1_tx_valid  <= 1'b1;
      while (!ep1_tx_ready) @(posedge clk);
      @(posedge clk);
      ep1_tx_valid  <= 1'b0;
    end
  endtask

  initial begin
    ep0_tx_valid = 1'b0; ep1_tx_valid = 1'b0;
    ep0_tx_data = 32'h0; ep1_tx_data = 32'h0;
    ep0_tx_dest = '0; ep1_tx_dest = '0;

    wait (rst_n);
    repeat (5) @(posedge clk);

    // Send multiple flits to ep0 to overflow and trigger Must‑Sink
    send_ep1(16'h1100, 32'h1111_0001);
    send_ep1(16'h1100, 32'h1111_0002);
    send_ep1(16'h1100, 32'h1111_0003);
    send_ep1(16'h1100, 32'h1111_0004);

    begin
      int tcnt;
      tcnt = 0;
      while (!ep0_rx_err && (tcnt < 200)) begin
        @(posedge clk);
        tcnt++;
      end
      if (!ep0_rx_err) $fatal("[TB] expected ep0_rx_err due to Must‑Sink drop");
    end

    $display("[TB] AXI‑MailboxFabric Must‑Sink test complete");
    $finish;
  end

endmodule
